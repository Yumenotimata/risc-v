module Decoder();
endmodule