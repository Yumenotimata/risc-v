module Execute();
endmodule