module Alu();
endmodule