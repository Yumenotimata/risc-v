module Fetch();
endmodule