`timescale 1ns/1ps
`include "core.v"
  
module startup;

    parameter step = 10;
    parameter ticks = 5000;
    parameter memory_hex = "build/riscv-tests-hex/rv32ui-p-sll.hex";
    parameter result_file_path = "result/rv32ui-p-sll.txt";

    reg clk;
    reg rst;

    Core core(
        .clk(clk),
        .rst(rst)
        );
    initial begin
        $readmemh(memory_hex,core.memory.m,16'h0,16'hffff);
    end

    integer i;
    initial
        begin
            $dumpfile("vcd/rv32ui-p-sll.vcd");
            $dumpvars(0,core);
            for(i=0;i<32;i++) begin
               $dumpvars(1,core.memory.m[i]);
            end
            for(i=0;i<31;i++) begin
                $dumpvars(2,core.rs[i]);
            end
            for(i=0;i<31;i++) begin
            //    $dumpvars(3,core.csr[i]);
            end
            $dumpvars(3,core.csr[12'h305]);
            $dumpvars(4,core.csr[305]);
        end

    initial
        begin
            clk = 1'b1;
            forever
                begin
                    #(step/2) clk = !clk;
                end
        end

    initial
        begin
            rst = 1'b0;
            repeat (1) @(posedge clk) rst <= 1'b1;
            @(posedge clk) rst <= 1'b0;
        end

    integer fp;

    initial
       begin
            repeat (ticks) @(posedge clk);
            fp = $fopen(result_file_path);
            if(core.rs[3] == 32'b1) begin
                $fdisplay(fp,"passed");
            end else begin
                $fdisplay(fp,"failed");
            end
            $finish();
            $fclose(fp);
        end

endmodule