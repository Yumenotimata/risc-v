module MemoryAccess();
endmodule