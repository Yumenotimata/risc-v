module MemoryAccess();

    wire [31:0] 

endmodule