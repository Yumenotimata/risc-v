module Decoder(
    input wire decoder_valid,
    input reg [31:0] decode_instruction
);

    always @(posedge decoder_valid) begin
        
    end

endmodule