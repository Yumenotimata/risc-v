module WriteBack();
endmodule